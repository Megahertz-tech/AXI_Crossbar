/// AXI Error Slave
///
/// This module always responds with an AXI error for transactions that are sent to it.
/// It's used to handle decode errors and invalid connections in the crossbar.
/// The module accepts transactions and immediately responds with decode errors.
///
/// Features:
/// - Configurable error response type
/// - Support for atomic operations (ATOPs)
/// - Configurable response data pattern
/// - Flow control to prevent resource exhaustion
///
/// TODO: Students should complete the implementation to properly handle
/// all AXI transactions and generate appropriate error responses.

module axi_err_slv #(
  parameter int unsigned          AxiIdWidth  = 0,                    // AXI ID Width
  parameter type                  axi_req_t   = logic,                // AXI 4 request struct, with atop field
  parameter type                  axi_resp_t  = logic,                // AXI 4 response struct
  parameter axi_pkg::resp_t       Resp        = axi_pkg::RESP_DECERR, // Error generated by this slave.
  parameter int unsigned          RespWidth   = 32'd64,               // Data response width, gets zero extended or truncated to r.data.
  parameter logic [RespWidth-1:0] RespData    = 64'hCA11AB1EBADCAB1E, // Hexvalue for data return value
  parameter bit                   ATOPs       = 1'b1,                 // Activate support for ATOPs.
  parameter int unsigned          MaxTrans    = 1                     // Maximum # of accepted transactions before stalling
) (
  input  logic      clk_i,   // Clock
  input  logic      rst_ni,  // Asynchronous reset active low
  input  logic      test_i,  // Testmode enable
  // slave port
  input  axi_req_t  slv_req_i,
  output axi_resp_t slv_resp_o
);

  // TODO: Define internal types
  typedef logic [AxiIdWidth-1:0] id_t;
  typedef struct packed {
    id_t           id;
    axi_pkg::len_t len;
  } r_data_t;

  // TODO: Handle ATOP filter if needed
  axi_req_t   err_req;
  axi_resp_t  err_resp;

  if (ATOPs) begin : gen_atop_filter
    // TODO: Students should implement ATOP filtering
    // For now, simple pass-through (students must enhance)
    axi_atop_filter #(
      .AxiIdWidth       ( AxiIdWidth  ),
      .AxiMaxWriteTxns  ( MaxTrans    ),
      .axi_req_t        ( axi_req_t   ),
      .axi_resp_t       ( axi_resp_t  )
    ) i_atop_filter (
      .clk_i,
      .rst_ni,
      .slv_req_i  ( slv_req_i   ),
      .slv_resp_o ( slv_resp_o  ),
      .mst_req_o  ( err_req     ),
      .mst_resp_i ( err_resp    )
    );
  end else begin : gen_no_atop
    assign err_req    = slv_req_i;
    assign slv_resp_o = err_resp;
  end

  // TODO: Implement FIFO structures for transaction tracking
  // W channel tracking
  logic    w_fifo_full, w_fifo_empty;
  logic    w_fifo_push, w_fifo_pop;
  id_t     w_fifo_data;

  // B channel tracking
  logic    b_fifo_full, b_fifo_empty;
  logic    b_fifo_push, b_fifo_pop;
  id_t     b_fifo_data;

  // R channel tracking
  r_data_t r_fifo_inp;
  logic    r_fifo_full, r_fifo_empty;
  logic    r_fifo_push, r_fifo_pop;
  r_data_t r_fifo_data;

  // R beat counter
  logic    r_cnt_clear, r_cnt_en, r_cnt_load;
  axi_pkg::len_t r_current_beat;
  logic    r_cnt_last;

  // TODO: Implement FIFO instances for transaction tracking
  fifo_v3 #(
    .DEPTH ( MaxTrans ),
    .dtype ( id_t     )
  ) i_w_fifo (
    .clk_i,
    .rst_ni,
    .flush_i    ( 1'b0       ),
    .testmode_i ( test_i     ),
    .full_o     ( w_fifo_full  ),
    .empty_o    ( w_fifo_empty ),
    .usage_o    (            ),
    .data_i     ( err_req.aw.id ),
    .push_i     ( w_fifo_push  ),
    .data_o     ( w_fifo_data  ),
    .pop_i      ( w_fifo_pop   )
  );

  fifo_v3 #(
    .DEPTH ( MaxTrans ),
    .dtype ( id_t     )
  ) i_b_fifo (
    .clk_i,
    .rst_ni,
    .flush_i    ( 1'b0       ),
    .testmode_i ( test_i     ),
    .full_o     ( b_fifo_full  ),
    .empty_o    ( b_fifo_empty ),
    .usage_o    (            ),
    .data_i     ( w_fifo_data  ),
    .push_i     ( b_fifo_push  ),
    .data_o     ( b_fifo_data  ),
    .pop_i      ( b_fifo_pop   )
  );

  fifo_v3 #(
    .DEPTH ( MaxTrans ),
    .dtype ( r_data_t )
  ) i_r_fifo (
    .clk_i,
    .rst_ni,
    .flush_i    ( 1'b0       ),
    .testmode_i ( test_i     ),
    .full_o     ( r_fifo_full  ),
    .empty_o    ( r_fifo_empty ),
    .usage_o    (            ),
    .data_i     ( r_fifo_inp   ),
    .push_i     ( r_fifo_push  ),
    .data_o     ( r_fifo_data  ),
    .pop_i      ( r_fifo_pop   )
  );

  // TODO: Implement beat counter for read responses
  counter #(
    .WIDTH     ( $bits(axi_pkg::len_t) ),
    .STICKY_EN ( 1'b0                  )
  ) i_r_cnt (
    .clk_i,
    .rst_ni,
    .clear_i ( r_cnt_clear      ),
    .en_i    ( r_cnt_en         ),
    .load_i  ( r_cnt_load       ),
    .down_i  ( 1'b0             ),
    .d_i     ( '0               ),
    .q_o     ( r_current_beat   ),
    .overflow_o ( /* unused */  )
  );

  // TODO: Implement error slave logic
  // Students need to implement:
  // 1. AW channel acceptance and W FIFO management
  // 2. AR channel acceptance and R FIFO management
  // 3. W channel consumption and B response generation
  // 4. R response generation with proper beat counting
  // 5. Error response generation with configurable response codes

  // PLACEHOLDER: Basic error response logic (students must enhance)
  always_comb begin
    // Default values
    err_resp = '0;
    w_fifo_push = 1'b0;
    w_fifo_pop = 1'b0;
    b_fifo_push = 1'b0;
    b_fifo_pop = 1'b0;
    r_fifo_push = 1'b0;
    r_fifo_pop = 1'b0;
    r_fifo_inp = '0;
    r_cnt_clear = 1'b0;
    r_cnt_en = 1'b0;
    r_cnt_load = 1'b0;

    // TODO: Students must implement complete error slave logic here
    // This is just a placeholder to prevent compilation errors

    // Basic AW channel handling
    err_resp.aw_ready = !w_fifo_full;
    w_fifo_push = err_req.aw_valid && err_resp.aw_ready;

    // Basic W channel handling
    err_resp.w_ready = !w_fifo_empty;
    if (err_req.w_valid && err_resp.w_ready && err_req.w.last) begin
      w_fifo_pop = 1'b1;
      b_fifo_push = 1'b1;
    end

    // Basic B channel response
    err_resp.b_valid = !b_fifo_empty;
    err_resp.b.id = b_fifo_data;
    err_resp.b.resp = Resp;
    err_resp.b.user = '0;
    b_fifo_pop = err_resp.b_valid && err_req.b_ready;

    // Basic AR channel handling
    err_resp.ar_ready = !r_fifo_full;
    r_fifo_inp.id = err_req.ar.id;
    r_fifo_inp.len = err_req.ar.len;
    r_fifo_push = err_req.ar_valid && err_resp.ar_ready;

    // Basic R channel response
    err_resp.r_valid = !r_fifo_empty;
    err_resp.r.id = r_fifo_data.id;
    err_resp.r.data = RespData;
    err_resp.r.resp = Resp;
    err_resp.r.last = (r_current_beat == r_fifo_data.len);
    err_resp.r.user = '0;

    if (err_resp.r_valid && err_req.r_ready) begin
      if (err_resp.r.last) begin
        r_fifo_pop = 1'b1;
        r_cnt_clear = 1'b1;
      end else begin
        r_cnt_en = 1'b1;
      end
    end
  end

  assign r_cnt_last = (r_current_beat == r_fifo_data.len);

  // TODO: Add parameter validation assertions
  // pragma translate_off
  `ifndef VERILATOR
  `ifndef XSIM
  initial begin : check_params
    assert (AxiIdWidth > 0) else
      $fatal(1, "AXI ID width must be > 0");
    assert (MaxTrans > 0) else
      $fatal(1, "Maximum transactions must be > 0");
    assert (RespWidth > 0) else
      $fatal(1, "Response width must be > 0");
  end
  `endif
  `endif
  // pragma translate_on

endmodule