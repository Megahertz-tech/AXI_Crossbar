/* ***********************************************************
    document:       axi_macrodef.sv
    author:         Celine (He Zhao) 
    Date:           09/29/2025
    Description:    encapsulate common Macros defination to  
                    define AXI and AXI-Lite Channel and  
                    Request/Response Structs  
**************************************************************/



