/* ***********************************************************
    document:       axi_inf.sv
    author:         Celine (He Zhao) 
    Date:           09/29/2025
    Description:    AXI Interface Definitions  
**************************************************************/



