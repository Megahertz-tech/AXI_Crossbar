/* ***********************************************************
    document:       tb_axi_regular_cfg.sv
    author:         Celine (He Zhao) 
    Date:           10/03/2025
    Description:    The configuration for the Regular transactions 
**************************************************************/
`ifndef __TB_AXI_REGULAR_CFG_SV__
`define __TB_AXI_REGULAR_CFG_SV__







`endif 
