/* ***********************************************************
    document:       axi_xbar_wrapper.sv
    author:         Celine (He Zhao) 
    Date:           10/03/2025
    Description:    wrapper for connection between DUT and TB  
**************************************************************/
`ifndef __AXI_XBAR_WRAPPER_SV__
`define __AXI_XBAR_WRAPPER_SV__

`include "axi_typedef_pkg.svh"
`include "axi_inf.sv"
`include "axi_macro_assign.svh"
module axi_xbar_wrapper
#(
  parameter int unsigned                                    AXI_USER_WIDTH      =  0,
  parameter axi_typedef_pkg::xbar_cfg_t                     Cfg                 = '0,
  parameter bit                                             ATOPS               = 1'b1,
  parameter bit [Cfg.NoSlvPorts-1:0][Cfg.NoMstPorts-1:0]    CONNECTIVITY        = '1,
  parameter type                                            rule_t              = axi_pkg::xbar_rule_32_t,
  localparam int unsigned                                   MstPortsIdxWidth    =
        (Cfg.NoMstPorts == 32'd1) ? 32'd1 : unsigned'($clog2(Cfg.NoMstPorts))
) (
  input  logic                                                      clk_i,
  input  logic                                                      rst_ni,
  input  logic                                                      test_i,
  input  rule_t [Cfg.NoAddrRules-1:0]                               addr_map_i,
  input  logic  [Cfg.NoSlvPorts-1:0]                                en_default_mst_port_i,
  input  logic  [Cfg.NoSlvPorts-1:0][MstPortsIdxWidth-1:0]          default_mst_port_i,
  axi_inf                                                           slv_ports [Cfg.NoSlvPorts-1:0],
  axi_inf                                                           mst_ports [Cfg.NoMstPorts-1:0]
);

  // TODO: Implement type definitions for interface-based connections
  localparam int unsigned AxiIdWidthMstPorts = Cfg.AxiIdWidthSlvPorts + $clog2(Cfg.NoSlvPorts);

  typedef logic [AxiIdWidthMstPorts     -1:0] id_mst_t;
  typedef logic [Cfg.AxiIdWidthSlvPorts -1:0] id_slv_t;
  typedef logic [Cfg.AxiAddrWidth       -1:0] addr_t;
  typedef logic [Cfg.AxiDataWidth       -1:0] data_t;
  typedef logic [Cfg.AxiDataWidth/8     -1:0] strb_t;
  typedef logic [AXI_USER_WIDTH         -1:0] user_t;

  // TODO: Define AXI channel types using macros
  `AXI_TYPEDEF_AW_CHAN_T(mst_aw_chan_t, addr_t, id_mst_t, user_t)
  `AXI_TYPEDEF_AW_CHAN_T(slv_aw_chan_t, addr_t, id_slv_t, user_t)
  `AXI_TYPEDEF_W_CHAN_T(w_chan_t, data_t, strb_t, user_t)
  `AXI_TYPEDEF_B_CHAN_T(mst_b_chan_t, id_mst_t, user_t)
  `AXI_TYPEDEF_B_CHAN_T(slv_b_chan_t, id_slv_t, user_t)
  `AXI_TYPEDEF_AR_CHAN_T(mst_ar_chan_t, addr_t, id_mst_t, user_t)
  `AXI_TYPEDEF_AR_CHAN_T(slv_ar_chan_t, addr_t, id_slv_t, user_t)
  `AXI_TYPEDEF_R_CHAN_T(mst_r_chan_t, data_t, id_mst_t, user_t)
  `AXI_TYPEDEF_R_CHAN_T(slv_r_chan_t, data_t, id_slv_t, user_t)
  `AXI_TYPEDEF_REQ_T(mst_req_t, mst_aw_chan_t, w_chan_t, mst_ar_chan_t)
  `AXI_TYPEDEF_REQ_T(slv_req_t, slv_aw_chan_t, w_chan_t, slv_ar_chan_t)
  `AXI_TYPEDEF_RESP_T(mst_resp_t, mst_b_chan_t, mst_r_chan_t)
  `AXI_TYPEDEF_RESP_T(slv_resp_t, slv_b_chan_t, slv_r_chan_t)

  // TODO: Implement interface conversion logic
  mst_req_t   [Cfg.NoMstPorts-1:0]  mst_reqs;
  mst_resp_t  [Cfg.NoMstPorts-1:0]  mst_resps;
  slv_req_t   [Cfg.NoSlvPorts-1:0]  slv_reqs;
  slv_resp_t  [Cfg.NoSlvPorts-1:0]  slv_resps; 
    /*
  slv_req_t   [Cfg.NoMstPorts-1:0]  mst_reqs;
  slv_resp_t  [Cfg.NoMstPorts-1:0]  mst_resps;
  mst_req_t   [Cfg.NoSlvPorts-1:0]  slv_reqs;
  mst_resp_t  [Cfg.NoSlvPorts-1:0]  slv_resps;
  */

  // Convert from struct-based to interface-based connections

  for (genvar i = 0; i < Cfg.NoMstPorts; i++) begin : gen_assign_mst
    `AXI_ASSIGN_FROM_REQ(mst_ports[i], mst_reqs[i])
    //`AXI_ASSIGN_TO_REQ(mst_reqs[i], mst_ports[i])
    `AXI_ASSIGN_TO_RESP(mst_resps[i], mst_ports[i])
    //`AXI_ASSIGN_FROM_RESP(mst_ports[i], mst_resps[i])
  end
  for (genvar i = 0; i < Cfg.NoSlvPorts; i++) begin : gen_assign_slv
    `AXI_ASSIGN_TO_REQ(slv_reqs[i], slv_ports[i])
        //assign slv_ports[i].aw_ready = slv_resps[i].aw_ready;
        //assign slv_ports[i].w_ready = slv_resps[i].w_ready;
        //assign slv_ports[i].b_valid = slv_resps[i].b_valid;
        //assign slv_ports[i].b_id = slv_resps[i].b.id;
        //assign slv_ports[i].b_resp = slv_resps[i].b.resp;
        //assign slv_ports[i].b_user = slv_resps[i].b.user;
        //assign slv_ports[i].ar_ready = slv_resps[i].ar_ready;
        //assign slv_ports[i].r_valid = slv_resps[i].r_valid;
        //assign slv_ports[i].r_id = slv_resps[i].r.id;
        //assign slv_ports[i].r_data = slv_resps[i].r.data;
        //assign slv_ports[i].r_resp = slv_resps[i].r.resp;
        //assign slv_ports[i].r_last = slv_resps[i].r.last;
        //assign slv_ports[i].r_user = slv_resps[i].r.user;
    `AXI_ASSIGN_FROM_RESP(slv_ports[i], slv_resps[i])
    //`AXI_ASSIGN_TO_RESP(slv_resps[i], slv_ports[i])
  end

  // TODO: Instantiate the main crossbar
  //{{{ 
  axi_xbar #(
    .Cfg  (Cfg),
    .ATOPs          ( ATOPS         ),
    .Connectivity   ( CONNECTIVITY  ),
    .slv_aw_chan_t  ( slv_aw_chan_t ),
    .mst_aw_chan_t  ( mst_aw_chan_t ),
    .w_chan_t       ( w_chan_t      ),
    .slv_b_chan_t   ( slv_b_chan_t  ),
    .mst_b_chan_t   ( mst_b_chan_t  ),
    .slv_ar_chan_t  ( slv_ar_chan_t ),
    .mst_ar_chan_t  ( mst_ar_chan_t ),
    .slv_r_chan_t   ( slv_r_chan_t  ),
    .mst_r_chan_t   ( mst_r_chan_t  ),
    .slv_req_t      ( slv_req_t     ),
    .slv_resp_t     ( slv_resp_t    ),
    .mst_req_t      ( mst_req_t     ),
    .mst_resp_t     ( mst_resp_t    ),
    .rule_t         ( rule_t        )
  ) i_xbar (
    .clk_i,
    .rst_ni,
    .test_i,
    .slv_ports_req_i  (slv_reqs ),
    .slv_ports_resp_o (slv_resps),
    .mst_ports_req_o  (mst_reqs ),
    .mst_ports_resp_i (mst_resps),
    .addr_map_i,
    .en_default_mst_port_i,
    .default_mst_port_i
  );
  //}}}

endmodule 

`endif 
