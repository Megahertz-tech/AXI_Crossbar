/* ***********************************************************
    document:       tb_axi_cfg_base.sv
    author:         Celine (He Zhao) 
    Date:           10/03/2025
    Description:     
**************************************************************/
`ifndef __TB_AXI_CFG_BASE_SV__
`define __TB_AXI_CFG_BASE_SV__
`include "tb_axi_macro_define_pkg.svh"
class tb_axi_cfg_base extends uvm_object;
    `uvm_object_utils(tb_axi_cfg_base)
    
    ob_construct(tb_axi_cfg_base)

    
endclass 

`endif 
