/* ***********************************************************
    document:       .sv
    author:         Celine (He Zhao) 
    Date:           10/03/2025
    Description:     
**************************************************************/
`ifndef ____
`define 







`endif 
