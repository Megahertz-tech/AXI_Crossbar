/* ***********************************************************
    document:       axi_xbar_default_slave.sv
    author:         Celine (He Zhao) 
    Date:           10/03/2025
    Description:     
**************************************************************/
`ifndef __AXI_XBAR_DEFAULT_SLAVE_SV__
`define __AXI_XBAR_DEFAULT_SLAVE_SV__

module axi_xbar_default_slave #(
  parameter int unsigned          AxiIdWidth  = 0,                    // AXI ID Width
  parameter type                  axi_req_t   = logic,                // AXI 4 request struct, with atop field
  parameter type                  axi_resp_t  = logic,                // AXI 4 response struct
  parameter axi_pkg::resp_t       Resp        = axi_pkg::RESP_DECERR, // Error generated by this slave.
  parameter int unsigned          RespWidth   = 32'd64,               // Data response width, gets zero extended or truncated to r.data.
  parameter logic [RespWidth-1:0] RespData    = 64'hCA11AB1EBADCAB1E, // Hexvalue for data return value
  //parameter bit                   ATOPs       = 1'b1,                 // Activate support for ATOPs.
  parameter int unsigned          MaxTrans    = 1                     // Maximum # of accepted transactions before stalling
) (
  input  logic      clk_i,   // Clock
  input  logic      rst_ni,  // Asynchronous reset active low
  input  logic      test_i,  // Testmode enable
  // slave port
  input  axi_req_t  slv_req_i,
  output axi_resp_t slv_resp_o
);

    typedef logic [AxiIdWidth-1:0] id_t;
    typedef struct packed {
        id_t                id;
        axi_pkg::len_t      len;
    } r_data_t;

    axi_req_t   err_req;

    axi_atomic_filter #(
        .axi_req_t          ( axi_req_t   )
    ) i_atomic_filter (
        .clk_i,
        .rst_ni,
        .slv_req_i          ( slv_req_i   ),
        .filtered_req_o     ( err_req     )
    );

    //{{{ pseudo code
    /*  non atomic aw:                          
            aw_id: for b 
        ar: 
            ar_id, ar_len for r 
        atomic aw: 
            aw_id: for b        (atomic store)
            aw_id, aw_len for r (atomic load, swap, compare)
            
        so: axi_atop_filter do the job as following 
              aw: 
                | if(is non-atomic || is atomic-store)
                |      do nothing.
                | else 
                |      assign req_i.ar_id  = req_i.aw_id
                |      if(is atomic-compare)
                |        assign req_i.ar_len = req_i.aw_len >> 1  
                |      else 
                |        assign req_i.ar_len = req_i.aw_len
              ar: do nothing. 
        
        so: axi_xbar_default_slave module do jobs as following
             aw & w & b cooperate: 
                | w_fifo: depth:      MaxTrans    
                |         data type:  aw_id 
                |         push_en:    
                |         pop_en:     
                | b_fifo: depth:      MaxTrans
                |         data_type:  aw_id
                |         push_en:    
                |         pop_en:     
                | output: aw_ready, w_ready, b_valid, b_id, b_resp, b_user
             ar (both ar and aw atomic load, swap, compare) 
             ar & r cooerate: 
                | r_fifo: depth:      MaxTrans
                |         data_type:  {ar_id, ar_len}
                |         push_en:    
                |         pop_en:     
                | output: ar_ready, r_valid, r_id, r_data, r_last, r_resp, r_user
    */
    //}}}
    // AW state machine 
    // W state machine  
    // B state machine  
    // AR state machine 
    typedef enum logic[3:0] {
        AW_IDLE                     = 4'b0001, 
        AW_APPROVE                  = 4'b0010, // non-atomic aw
        AW_ATOP_STORE_APPROVE       = 4'b0100, // atomic aw store
        AW_ATOP_NONE_STORE_APPROVE  = 4'b1000  // atomic aw load, swap, compare 
    } aw_state_e;
    typedef enum logic[2:0] {
        AR_IDLE                     = 3'b001,
        AR_APPROVE                  = 3'b010, // ar 
        AR_FALLTHOUGH_TO_R          = 3'b100  // for atomic aw: r response
    } ar_state_e;
    typedef enum logic[3:0] {
        W_IDLE                      = 4'b0001, 
        W_ONE_TR                    = 4'b0010, // w: len == 0
        W_MULTI_TR                  = 4'b0100, // w: len >  0
        W_FALLTHOUGH_TO_B           = 4'b1000  // for atomic aw: b response 
    } w_state_e;
    typedef enum logic[1:0] {
        B_IDLE                      = 2'b01,
        B_APPROVE                   = 2'b10   // b
    } b_state_e;
    typedef enum logic[3:0] {
        R_IDLE                      = 4'b0001, 
        R_APPROVE                   = 4'b0010, // r: initiate  
        R_PROCESS_ONE_TRANSFER      = 4'b0100, // r: len == 0
        R_PROCESS_MULTI_TRANSFER    = 4'b1000  // r: len >  0 
    } r_state_e;
    enum {AW_I_BIT = 0, AW_A_BIT = 1,   AW_ASA_BIT = 2, AW_ANSA_BIT = 3 } aw_state_bit_e;
    enum {AR_I_BIT = 0, AR_A_BIT = 1,   AR_FT_BIT  = 2                  } ar_state_bit_e;
    enum {W_I_BIT  = 0,  W_O_BIT = 1,   W_M_BIT    = 2, W_FT_BIT    = 3 } w_state_bit_e;
    enum {B_I_BIT  = 0,  B_A_BIT = 1                                    } b_state_bit_e;
    enum {R_I_BIT  = 0,  R_A_BIT = 1,   R_POT_BIT  = 2, R_PMT_BIT   = 3 } r_state_bit_e;
    
    aw_state_e      aw_sta_cur,     aw_sta_nxt;
    w_state_e       w_sta_cur,      w_sta_nxt;
    b_state_e       b_sta_cur,      b_sta_nxt;
    ar_state_e      ar_sta_cur,     ar_sta_nxt;
    r_state_e       r_sta_cur,      r_sta_nxt;
    //{{{ aw
    id_t            aw_id_cur,              aw_id_nxt;            //for w_fifo
    r_data_t        aw_atomic_r_data_cur,   aw_atomic_r_data_nxt; //for ar state machine
    always_ff @(posedge clk_i or negedge rst_ni) begin 
        if(!rst_ni) begin
            aw_sta_cur              <= AW_IDLE;
            aw_id_cur               <= '0;
            aw_atomic_r_data_cur    <= '0;
        end else begin
            aw_sta_cur              <= aw_sta_nxt;
            aw_id_cur               <= aw_id_nxt;
            aw_atomic_r_data_cur    <= aw_atomic_r_data_nxt;
        end
    end
    logic push_aw_id_to_w_fifo_en;   //for w_fifo
    logic w_fifo_empty, w_fifo_full; //for w_fifo
    logic b_fifo_empty, b_fifo_full; //for b_fifo
    logic r_fifo_empty, r_fifo_full; //for r_fifo
    always_comb begin
        aw_sta_nxt              = aw_sta_cur;
        aw_id_nxt               = aw_id_cur;
        push_aw_id_to_w_fifo_en = 1'b0;
        aw_atomic_r_data_nxt    = aw_atomic_r_data_cur;
        unique case(1'b1)
            aw_sta_cur[AW_I_BIT]: begin
                if(err_req.aw_valid) begin
                    if(err_req.aw.atop[5:4] == 2'b00  && (!w_fifo_full)) begin
                        aw_sta_nxt = AW_APPROVE;
                        aw_id_nxt  = err_req.aw.id;
                    end else if(w_fifo_empty && (!b_fifo_full) && (!err_req.w_valid))begin
                        if(err_req.aw.atop[5:4] == 2'b01) begin
                            aw_sta_nxt  = AW_ATOP_STORE_APPROVE;
                            aw_id_nxt   = err_req.aw.id;
                        end else begin
                            if(ar_sta_cur == AR_IDLE && (!r_fifo_full) && (!err_req.ar_valid)) begin
                                aw_sta_nxt                  = AW_ATOP_NONE_STORE_APPROVE;
                                aw_id_nxt                   = err_req.aw.id;
                                aw_atomic_r_data_nxt.id     = err_req.ar.id;
                                aw_atomic_r_data_nxt.len    = err_req.ar.len;
                            end
                        end
                    end
                end
            end
            aw_sta_cur[AW_A_BIT]: begin   // AW_APPROVE
                aw_sta_nxt              = AW_IDLE;
                push_aw_id_to_w_fifo_en = 1'b1;
            end
            aw_sta_cur[AW_ASA_BIT]: begin // AW_ATOP_STORE_APPROVE
                aw_sta_nxt              = AW_IDLE;
                push_aw_id_to_w_fifo_en = 1'b1;
            end
            aw_sta_cur[AW_ANSA_BIT]: begin //AW_ATOP_NONE_STORE_APPROVE
                aw_sta_nxt              = AW_IDLE;
                push_aw_id_to_w_fifo_en = 1'b1;
            end
            default: begin end
        endcase
    end
    //}}}
    //{{{ w
    //w_fifo 
    logic pop_w_fifo_en;             //to b
    id_t  b_id_from_w_fifo;          //to b
    fifo_v3 #(
        .FALL_THROUGH   (0       ),
        .DEPTH          (MaxTrans),
        .dtype          (id_t    )
    ) i_w_fifo (
        .clk_i,
        .rst_ni,
        .flush_i        (1'b0                   ),
        .testmode_i     (test_i                 ),
        .push_i         (push_aw_id_to_w_fifo_en),
        .data_i         (aw_id_cur              ),
        .pop_i          (pop_w_fifo_en          ),
        .data_o         (b_id_from_w_fifo       ),
        .full_o         (w_fifo_full            ),
        .empty_o        (w_fifo_empty           ),
        .usage_o        (/*not used*/           )
    );

    always_ff @(posedge clk_i or negedge rst_ni) begin 
        if(!rst_ni) begin
            w_sta_cur <= W_IDLE;
        end else begin
            w_sta_cur <= w_sta_nxt;
        end
    end
    always_comb begin
        w_sta_nxt = w_sta_cur;
        pop_w_fifo_en = 1'b0;
        unique case(1'b1)
            w_sta_cur[W_I_BIT]: begin // W_IDLE
                if(err_req.w_valid && (!w_fifo_empty) && (!b_fifo_full)) begin
                    if(err_req.w.last) begin
                        w_sta_nxt = W_ONE_TR;
                    end else begin
                        w_sta_nxt = W_MULTI_TR;
                    end 
                end
                if((aw_sta_cur == AW_ATOP_STORE_APPROVE) || (aw_sta_cur == AW_ATOP_NONE_STORE_APPROVE)) begin
                    w_sta_nxt = W_FALLTHOUGH_TO_B;
                end
            end
            w_sta_cur[W_O_BIT]: begin // W_ONE_TR
                w_sta_nxt       = W_IDLE;
                pop_w_fifo_en   = 1'b1;
            end
            w_sta_cur[W_M_BIT]: begin // W_MULTI_TR
                if(err_req.w.last)  begin
                    w_sta_nxt       = W_IDLE;
                    pop_w_fifo_en   = 1'b1;
                end
            end
            w_sta_cur[W_FT_BIT]: begin // W_FALLTHROUGH_TO_B
                w_sta_nxt       = W_IDLE;
                pop_w_fifo_en   = 1'b1;
            end
            default: begin end 
        endcase
    end 
    //}}}
    //{{{ b
    logic push_b_id_en;
    always_ff @(posedge clk_i or negedge rst_ni) begin 
        if(!rst_ni) begin
           push_b_id_en  <= 1'b0;
        end else begin
           push_b_id_en  <= pop_w_fifo_en;
        end
    end

    logic pop_b_id_en;
    id_t  b_id;
    fifo_v3 #(
        .FALL_THROUGH   (0          ),
        .DEPTH          (MaxTrans   ),
        .dtype          (id_t       )
    ) i_b_fifo (
        .clk_i,
        .rst_ni,
        .flush_i    (1'b0               ),
        .testmode_i (test_i             ),
        .push_i     (push_b_id_en       ),
        .data_i     (b_id_from_w_fifo   ), //from w_fifo 
        .pop_i      (pop_b_id_en        ), 
        .data_o     (b_id               ),
        .full_o     (b_fifo_full        ),
        .empty_o    (b_fifo_empty       ),
        .usage_o    (/*not used*/       )
    ); 
    always_ff @(posedge clk_i or negedge rst_ni) begin 
        if(!rst_ni) begin
            b_sta_cur <= B_IDLE;
        end else begin
            b_sta_cur <= b_sta_nxt;
        end
    end
    always_comb begin
        b_sta_nxt   = b_sta_cur;
        pop_b_id_en = 1'b0;
        unique case(1'b1) 
            b_sta_cur[B_I_BIT]: begin
                if(!b_fifo_empty) begin
                    b_sta_nxt   = B_APPROVE;
                    pop_b_id_en = 1'b1;
                end
            end
            b_sta_cur[B_A_BIT]: begin
                if(err_req.b_ready) begin
                    b_sta_nxt = B_IDLE;
                end
            end
            default: begin end 
        endcase
    end 
    //}}}
//{{{ ar
    r_data_t        r_data_cur,     r_data_nxt;
    always_ff @(posedge clk_i or negedge rst_ni) begin 
        if(!rst_ni) begin
            ar_sta_cur <= AR_IDLE;
            r_data_cur <= '0;
        end else begin
            ar_sta_cur <= ar_sta_nxt;
            r_data_cur <= r_data_nxt;
        end
    end
    logic   r_fifo_push_en;
    always_comb begin
        ar_sta_nxt      = ar_sta_cur;
        r_fifo_push_en  = 1'b0;
        r_data_nxt      = r_data_cur;
        unique case(1'b1)
            ar_sta_cur[AR_I_BIT]: begin // AR_IDLE
                if(err_req.ar_valid && (!r_fifo_full)) begin 
                    if(aw_sta_cur != AW_ATOP_NONE_STORE_APPROVE) begin
                        ar_sta_nxt      = AR_APPROVE;
                        r_data_nxt.id   = err_req.ar.id;
                        r_data_nxt.len  = err_req.ar.len;
                    end
                end
                if(aw_sta_cur == AW_ATOP_NONE_STORE_APPROVE) begin
                    ar_sta_nxt      = AR_FALLTHOUGH_TO_R;
                    r_data_nxt.id   = aw_atomic_r_data_cur.id;
                    r_data_nxt.len  = aw_atomic_r_data_cur.len;
                end
            end
            ar_sta_cur[AR_A_BIT]: begin // AR_APPROVE
                ar_sta_nxt      = AR_IDLE;
                r_fifo_push_en  = 1'b1;
            end
            ar_sta_cur[AR_FT_BIT]: begin// AR_FALLTHOUGH_TO_R
                ar_sta_nxt      = AR_IDLE;
                r_fifo_push_en  = 1'b1;
            end
            default: begin end 
        endcase
    end 
//}}}
    localparam int unsigned RLEN_WIDTH = $bits(axi_pkg::len_t) + 1;
//{{{ r 
    r_data_t    r_id_len;
    logic       r_pop_en;
    fifo_v3 #(
        .FALL_THROUGH   (0       ),
        .DEPTH          (MaxTrans),
        .dtype          (r_data_t)
    ) i_r_fifo (
        .clk_i,
        .rst_ni,
        .flush_i    (1'b0           ),
        .testmode_i (test_i         ),
        .push_i     (r_fifo_push_en ),
        .data_i     (r_data_cur     ), 
        .pop_i      (r_pop_en       ), 
        .data_o     (r_id_len       ),
        .full_o     (r_fifo_full    ),
        .empty_o    (r_fifo_empty   ),
        .usage_o    (/*not used*/   )
    );
    // transmit r
    /*      if(len = 0): one transfer  
            if(len > 0): multiple transfers 
    */
    always_ff @(posedge clk_i or negedge rst_ni) begin 
        if(!rst_ni) begin
            r_sta_cur <= R_IDLE;
        end else begin
            r_sta_cur <= r_sta_nxt;
        end
    end
    logic   r_last;
    always_comb begin
        r_sta_nxt = r_sta_cur;        
        r_pop_en  = 1'b0;
        unique case(1'b1)
            r_sta_cur[R_I_BIT]: begin // R_IDLE
                if(!r_fifo_empty) begin
                    r_sta_nxt = R_APPROVE;
                    r_pop_en  = 1'b1;
                end
            end
            r_sta_cur[R_A_BIT]: begin // R_APPROVE
                if(!r_id_len.len) begin
                    r_sta_nxt = R_PROCESS_ONE_TRANSFER;
                end
                else begin
                    r_sta_nxt = R_PROCESS_MULTI_TRANSFER;
                end
            end
            r_sta_cur[R_POT_BIT]: begin // R_PROCESS_ONE_TRANSFER
                if(err_req.r_ready) begin
                    r_sta_nxt = R_IDLE;
                end
            end
            r_sta_cur[R_PMT_BIT]: begin // R_PROCESS_MULTI_TRANSFER
                if(r_last) begin
                    r_sta_nxt = R_IDLE;
                end
            end
            default: begin end
        endcase
    end    
    logic [RLEN_WIDTH-1:0] r_length;
    always_ff @(posedge clk_i or negedge rst_ni) begin 
        if(!rst_ni) begin
            r_length    <= '0;
            r_last      <= 1'b0;
        end else if(r_sta_cur == R_PROCESS_MULTI_TRANSFER) begin
            if(err_req.r_ready) begin
                if(r_length == r_id_len.len) begin
                    r_last      <= 1'b1;
                    r_length    <= r_length + 1;
                end else if(r_length < r_id_len.len) begin
                    r_last      <= 1'b0;
                    r_length    <= r_length + 1;
                end
            end
        end else begin
            r_length    <= '0;
            r_last      <= 1'b0;
        end
    end
//}}}
    //output 
    always_comb begin
        slv_resp_o = '0;
        //aw_ready
        if(!(aw_sta_cur == AW_IDLE)) begin
            slv_resp_o.aw_ready = 1'b1;    
        end
        //w_ready
        if((w_sta_cur == W_ONE_TR) || (w_sta_cur == W_MULTI_TR)) begin
            slv_resp_o.w_ready = 1'b1;
        end
        //b_valid, b_id, b_resp, b_user
        if(b_sta_cur == B_APPROVE) begin
            slv_resp_o.b_valid  = 1'b1;
            slv_resp_o.b.id     = b_id;
            slv_resp_o.b.resp   = Resp;
            //b_user : by default
        end
        //ar_ready 
        if(ar_sta_cur == AR_APPROVE) begin
            slv_resp_o.ar_ready = 1'b1;
        end
        //r_valid, r_id, r_data, r_last, r_resp, r_user
        if(r_sta_cur == R_PROCESS_ONE_TRANSFER) begin
            slv_resp_o.r_valid  = 1'b1;
            slv_resp_o.r.id     = r_id_len.id;
            slv_resp_o.r.data   = RespData;
            slv_resp_o.r.last   = 1'b1;
            slv_resp_o.r.resp   = Resp;
            //r_user : by default
        end else if(r_sta_cur == R_PROCESS_MULTI_TRANSFER) begin
            slv_resp_o.r_valid  = 1'b1;
            slv_resp_o.r.id     = r_id_len.id;
            slv_resp_o.r.data   = RespData;
            slv_resp_o.r.last   = r_last;
            slv_resp_o.r.resp   = Resp;
            //r_user : by default
        end
    end




endmodule

`endif 
